
module floatingPoint_tb();
reg [15:0]a,b;
reg clk,op;
wire [15:0]s;

floatingPoint fp(a,b,op,s,clk);

initial begin
op=1'b0;
a=16'b0100101100100100; //exp more man more 
b=16'b0100011011001100; //a+b=0100110101000101; a-b=0100011101111100; -a+b= 1100011101111100; -a-b=1100110101000101
//op=1'b1;
#5
a=16'b0100100100100100; //exp more man less 
b=16'b0100011011001100; //a+b=0100110001000101; a-b=0100001011111000; -a+b= 1100001011111000; -a-b=1100110001000101
//op=1'b1;
#5
a=16'b0100011100100100; //exp less man more 
b=16'b0100101011001100; //a+b=0100110100101111; a-b=1100011001110100; -a+b= 0100011001110100; -a-b=1100110100101111
//op=1'b1;
#5
a=16'b0100010100100100; //exp less man less 
b=16'b0100101011001100; //a+b=0100110010101111; a-b=1011011101000000; -a+b= 0011011101000000; -a-b=1100110010101111
//op=1'b0;
#5
a=16'b0100011100100100; //exp equal man more 
b=16'b0100011011001100; //a+b=0100101011111000; a-b=0011010110000000; -a+b= 1011010110000000; -a-b=1100101011111000
//op=1'b0;
#5
a=16'b0100010100100100; //exp equal man less 
b=16'b0100011011001100; //a+b=0100100111111000; a-b=1011111010100000; -a+b= 0011111010100000; -a-b=1100100111111000
#5
a=16'b0100101100100100; //exp more man becomes equal when we shift
b=16'b0100011001001000; 
#5
a=16'b0100011100100100; //exp equal man equal 
b=16'b0100011100100100; //a+b=0100101100100100; a-b=0000000000000000; -a+b= 1000000000000000; -a-b=1100101100100100
#5
a=16'b0111111100100100; // when exponent is 31 ->NaN 
b=16'b0100011100100100;
#5
a=16'b0111110000000000; // exp all 1, man all zeros-> infinity 
b=16'b0100011100100100;
#5
a=16'b0000000000000000; // exp all 0, man all zeros-> 0 
b=16'b0100011100100100;
end	

initial begin
clk=0;
#1 clk=~clk;

end

initial begin
$dumpfile("test1.vcd");
$dumpvars(0,floatingPoint_tb);
$monitor("time=%2d op=%b, a=%b, b=%b, s=%b",$time, op,a,b,s);
end

endmodule

